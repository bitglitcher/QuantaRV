
module core
(

);

regfile regfile_0
( 
    .clk(),
    .rd(),
    .rd_d(),
    .wr(),
    .rs1(),
    .rs2(),
    .rs1_d(),
    .rs2_d()
);



endmodule