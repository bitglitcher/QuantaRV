
`ifndef __DEBUG__PORT__SV__
`define __DEBUG__PORT__SV__

`ifndef ALTERA_RESERVED_QIS
    `define __sim__
    `define DEBUG_PORT
    `define MEMORY_DEBUG_MSGS
`endif

`endif